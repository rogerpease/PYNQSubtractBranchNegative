`ifndef SBNModule_tb_include_vh_
`define SBNModule_tb_include_vh_

//Configuration current bd names
`define BD_NAME SBNModule_bfm_1
`define BD_INST_NAME SBNModule_bfm_1_i
`define BD_WRAPPER SBNModule_bfm_1_wrapper

//Configuration address parameters
`endif
